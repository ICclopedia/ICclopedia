Transistors characterization NMOS transistor simulation testbench

.INCLUDE ./simulation_netlist.spice

* Interactive simulation main entry *
.CONTROL

* Make a directory for our output simulation files and switch to it
shell mkdir -p results 
cd results/
* Generic prefix for our output files
set generic_prefix = 'simulation'

echo 
echo '----'
echo 'DC analysis sweep: Normalized Id vs. Vds for different Vgs bias'
echo '----'
echo 

* Choose parameters to save: 
* first DC parameters (needs to be done prior to sims)
* then lumped AC capacitance parameters (to ground)
* then relative AC capacitance parameters among terminals
save all @m1[gm] @m1[gmbs] @m1[gds] @m1[id] @m1[vgs] @m1[vds] @m1[vbs] @m1[vth] @m1[vdsat]
+        @m1[cgg] @m1[cdd] @m1[css] @m1[cbb]
+        @m1[cgs] @m1[cgd] @m1[cgb]
+        @m1[cdg] @m1[cds] @m1[cdb]
+        @m1[csg] @m1[csd] @m1[csb]

let vds_start = 0
let vds_end = 1.3
let vds_increment = 0.05
let vds_length=((vds_end-vds_start)/vds_increment)+1

let vgs_start = 0.1
let vgs_end = 1.3
let vgs_increment = 0.1
let vgs_length=((vgs_end-vgs_start)/vgs_increment)+1

DC Vds $&vds_start $&vds_end $&vds_increment Vgs $&vgs_start $&vgs_end $&vgs_increment 
let vdsat = @m1[vdsat]
reshape vdsat [$&vgs_length][$&vds_length]
let ngvec = ng
reshape ngvec [$&vgs_length][$&vds_length]
let vth = @m1[vth]
reshape vth [$&vgs_length][$&vds_length]

echo 'Vdsat values for each Vgs'
echo 
let index = 0
while index < vgs_length
    let vgs_point=ngvec[index][26]
    let vdsat_point=vdsat[index][26]
    let vth_point=vth[index][26]
    let veff_point=vgs_point-vth_point
    echo "Vgs: At Vgs: $&vgs_point V, Vdsat(@Vds=Vdd): $&vdsat_point"
    echo
    let index=index+1
end

* Plotting normalized Ids vs Vgs for different Vgs traces
setscale nd ; set our plot scale (i.e. x axis to the nd vector)
setcs xlabel = 'Drain to Source Voltage (V)'
setcs ylabel = 'Normalized Drain Current (mA/um)'
setcs title = 'DC Analysis: Normalized Drain Current vs Drain to Source Voltage' 
set filename = {$generic_prefix}{'_dc_analysis'}
set gnuplot_terminal = 'eps'
gnuplot $filename (-Vds#branch*1e+03)/(@m1[w]*1e6) title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing DC transfer characteristics data to a textfile'
set filetype=ascii
set filename = {$generic_prefix}{'_dc_analysis.raw'}
write $filename

echo 
echo '----'
echo 'DC Analysis: Transistor parameters sweep vs. Vgs (for different Vbs)'
echo '----'
echo 

* Plot y vs xscale
set xscale="veff"
* General plotting properties for postcript printout
* Needed for printing versus arbitrary x-axis (gnuplot does not work)
set hcopydevtype=postscript
set hcopypscolor = 1 

let vgs_start = 0.05
let vgs_end = 1.3
let vgs_increment = 0.05
let vgs_length=((vgs_end-vgs_start)/vgs_increment)+1

let vbs_start = -1.3
let vbs_end = 0
let vbs_increment = 0.1
let vbs_length=abs((vbs_end-vbs_start)/vbs_increment)+1

DC Vgs $&vgs_start $&vgs_end $&vgs_increment Vbs $&vbs_start $&vbs_end $&vbs_increment 
$ Gather main device parameters
let vth=@m1[vth][vgs_length-1]
echo "Vth: $&vth V"

$ Calculate important design parameters afterwards
let veff=ng-@m1[vth]
let gmtot=@m1[gm]+@m1[gmbs]           ; must account for back-gate transconductance
let gmid=(gmtot)/@m1[id]
let gmw=(gmtot)/(@m1[w]*@m1[m]*1e6)   ; in um
let ao=20*log10(abs(gmtot/@m1[gds]))  ; in dB

$ Note these approximations only work in active-sat
let ft=gmtot/(2*pi*abs(@m1[cgg]))
let fc=1/(2*pi*(1/@m1[gds])*((abs(@m1[cdg]))+(abs(@m1[cds]))+(abs(@m1[cdb]))))
let fom=gmid*ft

echo 'Plotting transistor parameters sweep'
setscale $xscale
foreach parameter gmid gmw ao ft fc fom
    echo
    echo "Plotting $parameter vs $xscale"
    setcs xlabel = "$xscale"
    setcs ylabel = "$parameter"
    setcs title = "$parameter vs. $xscale"
    set filename = "{$generic_prefix}_{$parameter}_{vbs_analysis}"
    plot dc2.$parameter
    hardcopy $filename{.ps} dc2.$parameter
    +    title $title xlabel $xlabel ylabel $ylabel 
end

echo 
echo '----'
echo 'DC Analysis: Transistor parameters sweep vs. Vgs (for different lengths)'
echo '----'
echo 

let vgs_start = 0.05
let vgs_end = 1.3
let vgs_increment = 0.05
let vgs_length=((vgs_end-vgs_start)/vgs_increment)+1

* For each transistor length, sweep:
*   - vgs from 0.05 to 1.3V in 0.05v
* foreach m_l $&m_lsize
foreach m_l 130n 180n 250n 350n 500n 700n 1u 1.5u 2u 3u
    alter @M1[L] = $m_l
    DC Vgs $&vgs_start $&vgs_end $&vgs_increment 
    $ Gather main device parameters
    let vth=@m1[vth][vgs_length-1]
    echo "Vth: $&vth V"

    $ Calculate important design parameters afterwards
    let veff=ng-@m1[vth]
    let gmid=@m1[gm]/@m1[id]
    let gmw=@m1[gm]/@m1[w]
    let ao=20*log10(@m1[gm]/@m1[gds])   ;in dB
    $ Note these approximations only work in active-sat
    $ put in log form 
    let ft=log10(@m1[gm]/(2*pi*abs(@m1[cgg])))
    let fc=log10(1/(2*pi*(1/@m1[gds])*((abs(@m1[cdg]))+(abs(@m1[cds]))+(abs(@m1[cdb])))))
    let fom=log10(gmid*ft)
    $ Update secscale for the current plot
    setscale $xscale
end

foreach parameter gmid ao ft fc fom
    echo "Plotting $parameter vs $xscale"
    setcs xlabel = "$xscale"
    setcs ylabel = "$parameter"
    setcs title = "$parameter vs. $xscale"
    set filename = "{$generic_prefix}_{$parameter}_{length_analysis}"
    echo $filename
    set multiple_plots="dc3.$parameter dc4.$parameter dc5.$parameter dc6.$parameter dc7.$parameter dc8.$parameter dc9.$parameter dc10.$parameter dc11.$parameter dc12.$parameter"
    plot $multiple_plots 
    hardcopy $filename{.ps} $multiple_plots 
    +    title $title xlabel $xlabel ylabel $ylabel 
end

echo '* Writing all simulation data to a textfile'
set filetype=ascii
set filename = {$generic_prefix}{'_transistor_parameters.raw'}
write $filename
* back to main directory
cd ../

.ENDC
