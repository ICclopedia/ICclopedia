* IC Resistor model and parameters 
* From: Designing Analog Chips by Hans Camenzind. 
* Reference: http://www.designinganalogchips.com/

* 3 Section/segment lumped model for integrated resistor 
.SUBCKT rcv 1 2
* dev   <nets>  model   expr
* --------------------------
R1      1 4     rb      {m/3}
R2      4 5     rb      {m/3}
R3      5 6     rb      {m/3}
V1      6 2 0
B1      6 1     i=i(v1)*(0.0033*((v(3)-(v(1)+v(2))/2))^0.6)
D1      1 3     drsub   {m/2}
D2      4 3     drsub   {m}
D3      5 3     drsub   {m}
D4      6 3     drsub   {m/2}
.ENDS

.MODEL drsub D is=1e-16 rs=50 cjo=2.7e-14 m=0.38 vj=0.6

