* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  /n_pos /0 1.3V		
I1  /n_pos /n1 50uA		
V2  /n2 /0 1.3V		
M1  /n1 /n1 /0 /0 L=5U W=2U		;Node Sequence Spec.<d,g,s,b>
M2  /n2 /n1 /0 /0 L=5U W=2U		;Node Sequence Spec.<d,g,s,b>

.end
