* Lateral PNP Wilson Current Mirror SPICE Netlist

.INCLUDE ../device_parameter_libraries/bipolar_20v_process.spice

* Circuit Elements: Devices
* dev <nets>               <values>
* ---------------------------------
V1    n_pos 0              5V		
I1    n3    0              50uA		
XQ1   n1    n3 n1  n_pos 0 split_coll_lat_pnp1 
XQ2   n2    n3 n1  0       lat_pnp1
V2    n2    0              4V		

.END
