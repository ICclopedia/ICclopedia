* Source Degeneration Resistors Negative Feedback

.INCLUDE ../device_parameter_libraries/cmos_ptm_asu_130nm_tt.spice

* Circuit Elements: Devices
* dev <nets>        <values>
* --------------------------
I1    n_pos n1      50uA		
V1    n_pos 0       1.3V		
V2    n2    0       0.8225957V 
M1    n1    n1 n3 0 nmos w=5u l=2u 
M2    n2    n1 n4 0 nmos w=5u l=2u 
R1    n3    0       3kR
R2    n4    0       3kR

.END
