Simple MOS Current Mirror

.INCLUDE simple_mos_current_mirror_simulation_netlist.spice

* Interactive simulation main entry *
.CONTROL

* Make a directory for our output simulation files.
shell mkdir -p results 
* Generic prefix for our output files
set generic_prefix = 'results/simple_mos_current_mirror_simulation'

echo  '* Operating point analysis: Nominal current match '

OP                      
print all               

* Output current over constant input current (with matched vds load): should be 1 for best match.
print (v2#branch/v1#branch)

echo
echo '*Printing relevant transistor DC parameters table'
show m : gm,gmbs,gds,id,vgs,vds,vbs,vth,vdsat

echo 
echo '*Performing DC analysis sweep: Voltage dependence of current mirror'

DC V2 0V 1.3V 0.05V          ; Sweep Drain voltage from 0v to 1.3v in 0.05v increments.

* set our plot scale (i.e. x axis to the n2 vector)
setscale n2 
* plotting properties
set title = 'DC Analysis: Current Output vs Drain Voltage' 
set xlabel = 'Drain Voltage (V)'
set ylabel = 'Current Output (uA)'
set yhigh = 46
set ylow = 52
set filename = {$generic_prefix}{'_dc_analysis'}
set gnuplot_terminal = 'eps'

gnuplot $filename (v2#branch*-1e+06) ylimit $ylow $yhigh title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing all simulation data to a textfile'

set filetype=ascii
set filename = {$generic_prefix}{'_results.raw'}
write $filename

.ENDC
