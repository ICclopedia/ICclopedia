Transistors characterization NMOS transistor simulation testbench

.INCLUDE ./simulation_netlist.spice

* Interactive simulation main entry *
.CONTROL

* Make a directory for our output simulation files and switch to it
shell mkdir -p results 
cd results/
* Generic prefix for our output files
set generic_prefix = 'simulation'

echo '----'
echo '*Performing DC analysis sweep: Normalized Id vs. Vds for different Vgs bias'
echo '----'
let vds_start = 0
let vds_end = 1.3
let vds_increment = 0.05
let vds_length=((vds_end-vds_start)/vds_increment)+1

let vgs_start = 0.1
let vgs_end = 1.3
let vgs_increment = 0.1
let vgs_length=((vgs_end-vgs_start)/vgs_increment)+1

save all @m1[vdsat] @m1[vth]
DC Vds $&vds_start $&vds_end $&vds_increment Vgs $&vgs_start $&vgs_end $&vgs_increment 
let vdsat = @m1[vdsat]
reshape vdsat [$&vgs_length][$&vds_length]
let ngvec = ng
reshape ngvec [$&vgs_length][$&vds_length]
let vth = @m1[vth]
reshape vth [$&vgs_length][$&vds_length]

echo 'Vdsat values for each Vgs'
echo 
let index = 0
while index < vgs_length
    let vgs_point=ngvec[index][26]
    let vdsat_point=vdsat[index][26]
    let vth_point=vth[index][26]
    let veff_point=vgs_point-vth_point
    echo "Vgs: At Vgs: $&vgs_point V, Vdsat(@Vds=Vdd): $&vdsat_point"
    echo
    let index=index+1
end

* Plotting normalized Ids vs Vgs for different Vgs traces
setscale nd ; set our plot scale (i.e. x axis to the nd vector)
setcs xlabel = 'Drain to Source Voltage (V)'
setcs ylabel = 'Normalized Drain Current (mA/um)'
setcs title = 'DC Analysis: Normalized Drain Current vs Drain to Source Voltage' 
set filename = {$generic_prefix}{'_dc_analysis'}
set gnuplot_terminal = 'eps'
gnuplot $filename (-Vds#branch*1e+03)/(@m1[w]*1e6) title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing DC transfer characteristics data to a textfile'
set filetype=ascii
set filename = {$generic_prefix}{'_dc_analysis.raw'}
write $filename

echo '----'
echo '*Performing transistor parameters sweep: transistor parameters vs Vgs'
echo '----'

* Plot y vs xscale
set xscale="gmid"

let vgs_start = 0.05
let vgs_end = 1.3
let vgs_increment = 0.05
let vgs_length=((vgs_end-vgs_start)/vgs_increment)+1

* Store first DC parameters (needs to be done prior to sim)
* then lumped AC capacitance parameters (to ground)
* then relative AC capacitance parameters among terminals
save all @m1[gm] @m1[gmbs] @m1[gds] @m1[id] @m1[vgs] @m1[vds] @m1[vbs] @m1[vth] @m1[vdsat]
+        @m1[cgg] @m1[cdd] @m1[css] @m1[cbb]
+        @m1[cgs] @m1[cgd] @m1[cgb]
+        @m1[cdg] @m1[cds] @m1[cdb]
+        @m1[csg] @m1[csd] @m1[csb]

* For each transistor length, sweep:
*   - vgs from 0.05 to 1.3V in 0.05v
*foreach m_l $&m_lsize
foreach m_l 130n 180n 250n 350n 500n 700n 1u 1.5u 2u 3u
    alter @M1[L] = $m_l
    DC Vgs $&vgs_start $&vgs_end $&vgs_increment 
    $ Gather main device parameters
    let vth=@m1[vth][vgs_length-1]
    echo "Vth: $&vth V"
    let gm=@m1[gm]
    let id=@m1[id]
    let w=@m1[w]*1e6 ;in um
    let ro=1/@m1[gds]

    $ Calculate important design parameters afterwards
    let veff=ng-vth
    let gmid=gm/id
    let gmw=gm/w
    let ao=20*log10(gm*ro)   ;in dB
    $ Note these approximations only work in active-sat
    let ft=gm/(2*pi*abs(@m1[cgg]))
    let fc=1/(2*pi*ro*((abs(@m1[cdg]))+(abs(@m1[cds]))+(abs(@m1[cdb]))))
    let fom=gmid*ft
    $ Update secscale for the current plot
    setscale $xscale
end

* Plotting properties for postcript printout
* Needed for printing versus arbitrary x-axis (gnuplot does not work)
set hcopydevtype=postscript
set hcopypscolor = 1 

echo '----'
echo 'Performing transistor parameters sweep'
echo '----'
echo "Plotting gm/id vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'gm/Id transconductor current efficiency (S/A)' 
setcs title = "gm/Id vs. $xscale"
set filename = {$generic_prefix}{'_gmid_analysis'}
set multiple_plots="dc2.gmid dc3.gmid dc4.gmid dc5.gmid dc6.gmid dc7.gmid dc8.gmid dc9.gmid dc10.gmid dc11.gmid"
plot $multiple_plots
hardcopy $filename{.ps} $multiple_plots
+    title $title xlabel $xlabel ylabel $ylabel 

echo "Plotting gm/w vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'gm/W transconductor area efficiency (S/um)'
setcs title = "gm/W vs. $xscale"
set filename = {$generic_prefix}{'_gmw_analysis'}
set multiple_plots="dc2.gmw dc3.gmw dc4.gmw dc5.gmw dc6.gmw dc7.gmw dc8.gmw dc9.gmw dc10.gmw dc11.gmw"
plot $multiple_plots
hardcopy $filename{.ps} $multiple_plots
+    title $title xlabel $xlabel ylabel $ylabel 

echo "Plotting ao vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'ao transconductor intrinsic gain (dB)'
setcs title = "ao vs. $xscale"
set filename = {$generic_prefix}{'_ao_analysis'}
set multiple_plots="dc2.ao dc3.ao dc4.ao dc5.ao dc6.ao dc7.ao dc8.ao dc9.ao dc10.ao dc11.ao"
plot $multiple_plots
hardcopy $filename{.ps} $multiple_plots
+    title $title xlabel $xlabel ylabel $ylabel 

echo "Plotting Ft  vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'Ft transconductor intrinsic gain (MHz)'
setcs title = "Ft vs. $xscale"
set filename = {$generic_prefix}{'_ft_analysis'}
set multiple_plots="dc2.ft dc3.ft dc4.ft dc5.ft dc6.ft dc7.ft dc8.ft dc9.ft dc10.ft dc11.ft"
plot $multiple_plots ylog
hardcopy $filename{.ps} $multiple_plots ylog
+    title $title xlabel $xlabel ylabel $ylabel 


echo "Plotting Fc  vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'Fc transconductor intrinsic gain (MHz)'
setcs title = "Fc vs. $xscale"
set filename = {$generic_prefix}{'_fc_analysis'}
set multiple_plots="dc2.fc dc3.fc dc4.fc dc5.fc dc6.fc dc7.fc dc8.fc dc9.fc dc10.fc dc11.fc"
plot $multiple_plots ylog
hardcopy $filename{.ps} $multiple_plots ylog
+    title $title xlabel $xlabel ylabel $ylabel 

echo "Plotting FOM  vs $xscale"
setcs xlabel = "$xscale"
setcs ylabel = 'FOM: gmid x Ft' 
setcs title = "FOM vs. $xscale"
set filename = {$generic_prefix}{'_fom_analysis'}
set multiple_plots="dc2.fom dc3.fom dc4.fom dc5.fom dc6.fom dc7.fom dc8.fom dc9.fom dc10.fom dc11.fom"
plot $multiple_plots ylog 
hardcopy $filename{.ps} $multiple_plots ylog
+    title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing all simulation data to a textfile'
set filetype=ascii
set filename = {$generic_prefix}{'_transistor_parameters.raw'}
write $filename
* back to main directory
cd ../

.ENDC
