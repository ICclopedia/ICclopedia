* Simple PMOS Current Mirror

.INCLUDE ../device_parameter_libraries/cmos_ptm_asu_130nm_tt.spice

* Circuit Elements:  Devices
* dev <nets>         <values>
* --------------------------
V1    n_pos 0              1.3V		
I1    n1    0              50uA		
M1    n1    n1 n_pos n_pos pmos W=50u L=2u
M2    n2    n1 n_pos n_pos pmos W=50u L=2u
V2    n_pos n2             0.55957V

.END
