Lateral PNP Current Mirror

.INCLUDE lateral_pnp_current_mirror_simulation_netlist.spice

* Interactive simulation main entry *
.CONTROL

* Make a directory for our output simulation files.
shell mkdir -p results 
cd results

* Generic prefix for our output files
set generic_prefix = 'lateral_pnp_current_mirror_simulation'

echo  '* Operating point analysis: Current match '

OP                      
print all               

* Output current over constant input current (with 1V load): should be 1 for best match.
print (v2#branch/50e-06)

echo
echo '* DC analysis: Voltage dependence of current mirror'

DC V2 0V 4.89V 0.01V          ; Sweep Collector voltage from 0v to 5v in 0.01v increments.

* set our plot scale (i.e. x axis to the n2 vector)
setscale n2 
* plotting properties
setcs xlabel = 'Collector Voltage (V)'
setcs ylabel = 'Collector Current Output (uA)'
set xdel = 0.5
set yhigh = 60
set ylow = 41
set gnuplot_terminal = 'eps'

setcs title = 'DC Analysis: Collector Current Output vs Collector Voltage' 
set filename = {$generic_prefix}{'_dc_analysis_sweep'}
gnuplot $filename (v2#branch*1e+06) xdelta $xdel title $title xlabel $xlabel ylabel $ylabel 

setcs title = 'DC Analysis: Collector Current Output vs Collector Voltage (Zoom)' 
set filename = {$generic_prefix}{'_dc_analysis'}
gnuplot $filename (v2#branch*1e+06) ylimit $ylow $yhigh xdelta $xdel title $title xlabel $xlabel ylabel $ylabel 

echo '* Writing all simulation data to a textfile'

set filetype=ascii
set filename = {$generic_prefix}{'_results.raw'}
write $filename

.ENDC
