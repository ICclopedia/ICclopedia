* /media/camilo/data/workspaces/academia/self_study_courses/aic_1-analog_integrated_circuits/lab_assignments/3_current_mirrors/3_simple_mos_current_mirror/simple_mos_current_mirror.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu 14 Sep 2017 05:19:39 PM JST

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
V1  /n_pos /0 1.3V		
I1  /n_pos /n1 50uA		
V2  /n2 /0 1.3V		
M1  /n1 /n1 /0 /0 L=5U W=2U		;Node Sequence Spec.<d,g,s,b>
M2  /n2 /n1 /0 /0 L=5U W=2U		;Node Sequence Spec.<d,g,s,b>

.end
